`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company:       UPB
// Engineer:      Ovidiu Moldoveanu
//
// Create Date:   15:51:30 09/10/2021
// Design Name:   tester Baggage Drop
// Module Name:   tester
// Project Name:  Tema 1 - Baggage Drop
// Target Device: ISim
// Tool versions: 14.7
// Description:   tester for combinational module
////////////////////////////////////////////////////////////////////////////////

module adapter();

endmodule
